* SkyWater PDK
* Minimum size CMOS inverter
* VDD = 1.8 V, Lmin = 0.15um, Wn(min) = 0.42um

.lib /foss/pdks/sky130A/libs.tech/ngspice/sky130.lib.spice tt

*the voltage sources:
Vdd vdd gnd DC 1.8
V1 in gnd pulse(0 1.8 0p 20p 10p 1n 2n)

Xnot1 in vdd gnd inter not1
Xnot2 inter vdd gnd load not1

.subckt not1 A vdd vss y
xm02 y A vss vss sky130_fd_pr__nfet_01v8 l=0.15 w=0.42 as=0.126 ad=0.126 ps=1.44 pd=1.44
xm01 y A vdd vdd sky130_fd_pr__pfet_01v8 l=0.15 w=1.2 as=0.36 ad=0.36 ps=3 pd=3
.ends

* simulation command:
.tran 1ps 10ns 0 10p

.measure tran trise TRIG v(load) VAL={0.2*1.8} RISE=1 TARG v(load) VAL={0.8*1.8} RISE=1
.measure tran tfall TRIG v(load) VAL={0.8*1.8} FALL=1 TARG v(load) VAL={0.2*1.8} FALL=1
.measure tran tpHL  TRIG v(in)   VAL={0.5*1.8} FALL=1 TARG v(load) VAL={0.5*1.8} FALL=1
.measure tran tpLH  TRIG v(in)   VAL={0.5*1.8} RISE=1 TARG v(load) VAL={0.5*1.8} RISE=1
.measure tran tp_avg PARAM='(tpHL + tpLH)/2'

.control
run
plot in load

.endc
