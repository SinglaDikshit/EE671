magic
tech ihp-sg13g2
timestamp 1756313415
<< nwell >>
rect -96 -26 133 201
rect -96 -27 34 -26
<< pwell >>
rect -69 -49 33 -48
rect -69 -109 92 -49
rect -22 -111 92 -109
<< nmos >>
rect 30 -100 45 -58
<< pmos >>
rect 30 5 45 125
<< ndiff >>
rect -10 -65 30 -58
rect -10 -93 1 -65
rect 19 -93 30 -65
rect -10 -100 30 -93
rect 45 -65 85 -58
rect 45 -93 56 -65
rect 74 -93 85 -65
rect 45 -100 85 -93
<< pdiff >>
rect -10 117 30 125
rect -10 12 3 117
rect 19 12 30 117
rect -10 5 30 12
rect 45 45 85 125
rect 45 12 56 45
rect 72 12 85 45
rect 45 5 85 12
<< ndiffc >>
rect 1 -93 19 -65
rect 56 -93 74 -65
<< pdiffc >>
rect 3 12 19 117
rect 56 12 72 45
<< psubdiff >>
rect -50 -65 -10 -58
rect -50 -93 -39 -65
rect -21 -93 -10 -65
rect -50 -100 -10 -93
<< nsubdiff >>
rect -50 105 -10 125
rect -50 15 -40 105
rect -20 15 -10 105
rect -50 5 -10 15
<< psubdiffcont >>
rect -39 -93 -21 -65
<< nsubdiffcont >>
rect -40 15 -20 105
<< poly >>
rect 30 125 45 143
rect 30 -15 45 5
rect -5 -23 45 -15
rect -5 -39 2 -23
rect 22 -39 45 -23
rect -5 -46 45 -39
rect 30 -58 45 -46
rect 30 -120 45 -100
<< polycont >>
rect 2 -39 22 -23
<< metal1 >>
rect -27 148 103 151
rect -27 128 1 148
rect 22 128 61 148
rect 82 128 103 148
rect -27 127 103 128
rect -1 117 27 127
rect -1 107 3 117
rect -48 105 3 107
rect -48 15 -40 105
rect -20 15 3 105
rect -48 12 3 15
rect 19 12 27 117
rect -48 7 27 12
rect 49 45 77 50
rect 49 12 56 45
rect 72 12 77 45
rect -7 -23 30 -13
rect -7 -39 2 -23
rect 22 -39 30 -23
rect -7 -45 30 -39
rect 49 -58 77 12
rect -46 -63 -25 -60
rect -46 -65 28 -63
rect -46 -93 -41 -65
rect -21 -93 1 -65
rect 22 -93 28 -65
rect -46 -98 28 -93
rect 49 -65 81 -58
rect 49 -93 56 -65
rect 74 -93 81 -65
rect 49 -98 81 -93
rect -6 -117 28 -98
rect -24 -142 -1 -117
rect 19 -142 92 -117
rect -24 -143 92 -142
<< via1 >>
rect 1 128 22 148
rect 61 128 82 148
rect -41 -93 -39 -65
rect -39 -93 -21 -65
rect 1 -93 19 -65
rect 19 -93 22 -65
rect -1 -142 19 -117
<< metal2 >>
rect -28 148 103 153
rect -28 128 1 148
rect 22 128 61 148
rect 82 128 103 148
rect -28 127 103 128
rect -46 -65 29 -60
rect -46 -93 -41 -65
rect -21 -93 1 -65
rect 22 -93 29 -65
rect -32 -142 -1 -117
rect 19 -142 94 -117
rect -32 -149 94 -142
<< labels >>
flabel metal1 -5 -38 27 -23 0 FreeSans 80 0 0 0 A
port 1 nsew
flabel nwell -15 134 6 148 0 FreeSans 80 0 0 0 vdd
port 6 nsew
flabel metal2 -9 -136 17 -118 0 FreeSans 80 0 0 0 vss
port 7 nsew
flabel metal1 59 -40 69 -11 0 FreeSans 80 0 0 0 y
flabel metal1 59 -42 70 -15 0 FreeSans 80 0 0 0 y
port 8 nsew
<< end >>
