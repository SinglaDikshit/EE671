magic
tech ihp-sg13g2
timestamp 1756316239
<< poly >>
rect 91 125 128 132
rect 91 101 99 125
rect 123 124 128 125
rect 123 101 354 124
rect 91 94 128 101
<< polycont >>
rect 99 101 123 125
<< metal1 >>
rect 195 272 318 298
rect 91 125 128 132
rect 91 101 99 125
rect 123 101 128 125
rect 169 110 396 133
rect 91 99 128 101
rect 183 -6 319 27
<< metal2 >>
rect 195 272 318 298
rect 183 -6 319 27
use assgn2_trial  assgn2_trial_0 /foss/designs
timestamp 1756315725
transform 1 0 98 0 1 144
box -96 -149 133 201
use assgn2_trial  assgn2_trial_1
timestamp 1756315725
transform 1 0 326 0 1 145
box -96 -149 133 201
<< labels >>
flabel metal1 101 103 113 126 0 FreeSans 80 0 0 0 A
port 0 nsew
<< end >>
