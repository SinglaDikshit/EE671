* NGSPICE file created from str2.ext - technology: ihp-sg13g2

.subckt assgn2_trial vdd vss y a_n10_n92#
X0 y a_n10_n92# vss vss sg13_lv_nmos ad=0.11159p pd=0.93333u as=0.6315p ps=4.78u w=0.42u l=0.15u
**devattr s=6720,328 d=6720,328
X1 y a_n10_n92# vdd vdd sg13_lv_pmos ad=0.31881p pd=2.66667u as=1.118p ps=6.42u w=1.2u l=0.15u
**devattr s=19200,640 d=19200,640
C0 y a_n10_n92# 0.01838f
C1 vdd a_n10_n92# 0.10431f
C2 y vdd 0.12572f
C3 y vss 0.22148f
C4 vdd vss 0.22301f
C5 a_n10_n92# vss 0.27705f
.ends

.subckt str2 A
Xassgn2_trial_0 assgn2_trial_1/vdd VSUB assgn2_trial_1/y A assgn2_trial
Xassgn2_trial_1 assgn2_trial_1/vdd VSUB assgn2_trial_1/y A assgn2_trial
C0 assgn2_trial_1/y assgn2_trial_1/vdd 0.22759f
C1 assgn2_trial_1/vdd VSUB -0.03558f
C2 A assgn2_trial_1/vdd 0.15679f
C3 assgn2_trial_1/y VSUB 0.16698f
C4 A assgn2_trial_1/y 0.12528f
C5 A VSUB 0.08763f
C6 VSUB 0 0.02272f
C7 assgn2_trial_1/vdd 0 0.40157f
C8 assgn2_trial_1/y 0 0.38943f
C9 A 0 0.65227f
.ends

