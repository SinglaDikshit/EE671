* NGSPICE file created from str2.ext - technology: ihp-sg13g2

.subckt assgn2_trial vdd vss y a_n10_n92#
X0 y a_n10_n92# vss vss sg13_lv_nmos ad=0.11159p pd=0.93333u as=0.6315p ps=4.78u w=0.42u l=0.15u
**devattr s=6720,328 d=6720,328
X1 y a_n10_n92# vdd vdd sg13_lv_pmos ad=0.31881p pd=2.66667u as=1.118p ps=6.42u w=1.2u l=0.15u
**devattr s=19200,640 d=19200,640
.ends

.subckt str2 A
Xassgn2_trial_0 assgn2_trial_1/vdd VSUB assgn2_trial_1/y A assgn2_trial
Xassgn2_trial_1 assgn2_trial_1/vdd VSUB assgn2_trial_1/y A assgn2_trial
.ends

